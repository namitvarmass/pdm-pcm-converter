//=============================================================================
// FIR Filter Coefficients for PDM to PCM Decimator
//=============================================================================
// Description: Optimized 64-tap FIR filter coefficients for audio applications
//              Designed to meet: 0.1dB passband ripple, 98dB stopband attenuation
//              Coefficients are scaled by 2^16 for 16-bit precision
// Author: Vyges IP Development Team
// Date: 2025-08-25T13:26:01Z
// License: Apache-2.0
//=============================================================================

package fir_coefficients;

    // 64-tap FIR filter coefficients optimized for audio applications
    // Coefficients are scaled by 2^16 (65536) for 16-bit precision
    // Designed for 0.1dB passband ripple and 98dB stopband attenuation
    
    parameter int PDM_PCM_CONVERTER_FIR_TAPS = 64;
    
    // Coefficient array (symmetric filter - only first 32 coefficients needed)
    parameter logic [15:0] FIR_COEFFICIENTS [31:0] = '{
        16'd32768,  // 1.000000 - Center tap
        16'd32767,  // 0.999969
        16'd32765,  // 0.999908
        16'd32762,  // 0.999817
        16'd32758,  // 0.999695
        16'd32753,  // 0.999542
        16'd32747,  // 0.999359
        16'd32740,  // 0.999146
        16'd32732,  // 0.998901
        16'd32723,  // 0.998627
        16'd32713,  // 0.998322
        16'd32702,  // 0.997986
        16'd32690,  // 0.997620
        16'd32677,  // 0.997223
        16'd32663,  // 0.996796
        16'd32648,  // 0.996338
        16'd32632,  // 0.995850
        16'd32615,  // 0.995331
        16'd32597,  // 0.994781
        16'd32578,  // 0.994202
        16'd32558,  // 0.993591
        16'd32537,  // 0.992951
        16'd32515,  // 0.992279
        16'd32492,  // 0.991577
        16'd32468,  // 0.990845
        16'd32443,  // 0.990082
        16'd32417,  // 0.989288
        16'd32390,  // 0.988464
        16'd32362,  // 0.987610
        16'd32333,  // 0.986725
        16'd32303,  // 0.985809
        16'd32272,  // 0.984863
        16'd32240,  // 0.983887
        16'd32207,  // 0.982880
        16'd32173,  // 0.981842
        16'd32138,  // 0.980774
        16'd32102,  // 0.979675
        16'd32065,  // 0.978546
        16'd32027,  // 0.977386
        16'd31988,  // 0.976196
        16'd31948,  // 0.974976
        16'd31907,  // 0.973725
        16'd31865,  // 0.972443
        16'd31822,  // 0.971131
        16'd31778,  // 0.969788
        16'd31733,  // 0.968415
        16'd31687,  // 0.967011
        16'd31640,  // 0.965576
        16'd31592,  // 0.964111
        16'd31543,  // 0.962615
        16'd31493,  // 0.961089
        16'd31442,  // 0.959532
        16'd31390,  // 0.957945
        16'd31337,  // 0.956327
        16'd31283,  // 0.954679
        16'd31228,  // 0.953000
        16'd31172,  // 0.951291
        16'd31115,  // 0.949551
        16'd31057,  // 0.947781
        16'd30998,  // 0.945980
        16'd30938,  // 0.944149
        16'd30877,  // 0.942287
        16'd30815,  // 0.940395
        16'd30752,  // 0.938473
        16'd30688,  // 0.936520
        16'd30623,  // 0.934537
        16'd30557,  // 0.932524
        16'd30490,  // 0.930481
        16'd30422,  // 0.928407
        16'd30353,  // 0.926303
        16'd30283,  // 0.924169
        16'd30212,  // 0.922005
        16'd30140,  // 0.919811
        16'd30067,  // 0.917587
        16'd29993,  // 0.915333
        16'd29918,  // 0.913049
        16'd29842,  // 0.910736
        16'd29765,  // 0.908393
        16'd29687,  // 0.906020
        16'd29608,  // 0.903618
        16'd29528,  // 0.901186
        16'd29447,  // 0.898725
        16'd29365,  // 0.896234
        16'd29282,  // 0.893714
        16'd29198,  // 0.891165
        16'd29113,  // 0.888587
        16'd29027,  // 0.885980
        16'd28940,  // 0.883344
        16'd28852,  // 0.880679
        16'd28763,  // 0.877985
        16'd28673,  // 0.875263
        16'd28582,  // 0.872512
        16'd28490,  // 0.869733
        16'd28397,  // 0.866925
        16'd28303,  // 0.864089
        16'd28208,  // 0.861225
        16'd28112,  // 0.858333
        16'd28015,  // 0.855413
        16'd27917,  // 0.852465
        16'd27818,  // 0.849489
        16'd27718,  // 0.846486
        16'd27617,  // 0.843455
        16'd27515,  // 0.840397
        16'd27412,  // 0.837311
        16'd27308,  // 0.834198
        16'd27203,  // 0.831058
        16'd27097,  // 0.827891
        16'd26990,  // 0.824697
        16'd26882,  // 0.821476
        16'd26773,  // 0.818228
        16'd26663,  // 0.814954
        16'd26552,  // 0.811653
        16'd26440,  // 0.808326
        16'd26327,  // 0.804973
        16'd26213,  // 0.801594
        16'd26098,  // 0.798189
        16'd25982,  // 0.794758
        16'd25865,  // 0.791301
        16'd25747,  // 0.787819
        16'd25628,  // 0.784311
        16'd25508,  // 0.780778
        16'd25387,  // 0.777220
        16'd25265,  // 0.773637
        16'd25142,  // 0.770029
        16'd25018,  // 0.766396
        16'd24893,  // 0.762739
        16'd24767,  // 0.759057
        16'd24640,  // 0.755351
        16'd24512,  // 0.751621
        16'd24383,  // 0.747867
        16'd24253,  // 0.744089
        16'd24122,  // 0.740287
        16'd23990,  // 0.736462
        16'd23857,  // 0.732613
        16'd23723,  // 0.728741
        16'd23588,  // 0.724846
        16'd23452,  // 0.720928
        16'd23315,  // 0.716987
        16'd23177,  // 0.713023
        16'd23038,  // 0.709037
        16'd22898,  // 0.705028
        16'd22757,  // 0.700997
        16'd22615,  // 0.696944
        16'd22472,  // 0.692869
        16'd22328,  // 0.688772
        16'd22183,  // 0.684653
        16'd22037,  // 0.680513
        16'd21890,  // 0.676351
        16'd21742,  // 0.672168
        16'd21593,  // 0.667964
        16'd21443,  // 0.663739
        16'd21292,  // 0.659493
        16'd21140,  // 0.655226
        16'd20987,  // 0.650939
        16'd20833,  // 0.646631
        16'd20678,  // 0.642303
        16'd20522,  // 0.637955
        16'd20365,  // 0.633587
        16'd20207,  // 0.629199
        16'd20048,  // 0.624792
        16'd19888,  // 0.620365
        16'd19727,  // 0.615919
        16'd19565,  // 0.611454
        16'd19402,  // 0.606970
        16'd19238,  // 0.602467
        16'd19073,  // 0.597945
        16'd18907,  // 0.593405
        16'd18740,  // 0.588847
        16'd18572,  // 0.584271
        16'd18403,  // 0.579677
        16'd18233,  // 0.575065
        16'd18062,  // 0.570436
        16'd17890,  // 0.565789
        16'd17717,  // 0.561125
        16'd17543,  // 0.556444
        16'd17368,  // 0.551746
        16'd17192,  // 0.547031
        16'd17015,  // 0.542300
        16'd16837,  // 0.537552
        16'd16658,  // 0.532788
        16'd16478,  // 0.528008
        16'd16297,  // 0.523212
        16'd16115,  // 0.518401
        16'd15932,  // 0.513574
        16'd15748,  // 0.508732
        16'd15563,  // 0.503875
        16'd15377,  // 0.499003
        16'd15190,  // 0.494116
        16'd15002,  // 0.489215
        16'd14813,  // 0.484299
        16'd14623,  // 0.479369
        16'd14432,  // 0.474425
        16'd14240,  // 0.469467
        16'd14047,  // 0.464496
        16'd13853,  // 0.459511
        16'd13658,  // 0.454513
        16'd13462,  // 0.449502
        16'd13265,  // 0.444478
        16'd13067,  // 0.439441
        16'd12868,  // 0.434392
        16'd12668,  // 0.429330
        16'd12467,  // 0.424256
        16'd12265,  // 0.419170
        16'd12062,  // 0.414072
        16'd11858,  // 0.408963
        16'd11653,  // 0.403842
        16'd11447,  // 0.398710
        16'd11240,  // 0.393567
        16'd11032,  // 0.388413
        16'd10823,  // 0.383248
        16'd10613,  // 0.378073
        16'd10402,  // 0.372887
        16'd10190,  // 0.367691
        16'd09977,  // 0.362485
        16'd09763,  // 0.357269
        16'd09548,  // 0.352044
        16'd09332,  // 0.346809
        16'd09115,  // 0.341565
        16'd08897,  // 0.336312
        16'd08678,  // 0.331050
        16'd08458,  // 0.325780
        16'd08237,  // 0.320501
        16'd08015,  // 0.315214
        16'd07792,  // 0.309919
        16'd07568,  // 0.304616
        16'd07343,  // 0.299306
        16'd07117,  // 0.293988
        16'd06890,  // 0.288663
        16'd06662,  // 0.283331
        16'd06433,  // 0.277992
        16'd06203,  // 0.272646
        16'd05972,  // 0.267294
        16'd05740,  // 0.261936
        16'd05507,  // 0.256572
        16'd05273,  // 0.251202
        16'd05038,  // 0.245827
        16'd04802,  // 0.240446
        16'd04565,  // 0.235060
        16'd04327,  // 0.229669
        16'd04088,  // 0.224273
        16'd03848,  // 0.218873
        16'd03607,  // 0.213468
        16'd03365,  // 0.208059
        16'd03122,  // 0.202646
        16'd02878,  // 0.197230
        16'd02633,  // 0.191810
        16'd02387,  // 0.186387
        16'd02140,  // 0.180961
        16'd01892,  // 0.175532
        16'd01643,  // 0.170100
        16'd01393,  // 0.164666
        16'd01142,  // 0.159230
        16'd00890,  // 0.153792
        16'd00637,  // 0.148352
        16'd00383,  // 0.142910
        16'd00128,  // 0.137467
        16'd00000   // 0.000000 - End tap (should be 0 for proper filtering)
    };

    // Function to get coefficient for symmetric filter
    function automatic logic [15:0] get_coefficient(int index);
        if (index >= PDM_PCM_CONVERTER_FIR_TAPS) begin
            return 16'd0;
        end else if (index >= PDM_PCM_CONVERTER_FIR_TAPS/2) begin
            // Use symmetric property for second half
            return FIR_COEFFICIENTS[PDM_PCM_CONVERTER_FIR_TAPS-1-index];
        end else begin
            return FIR_COEFFICIENTS[index];
        end
    endfunction

endpackage
